module xadac #(
) (
    input logic clk_i,
    input logic rst_ni
);


endmodule
