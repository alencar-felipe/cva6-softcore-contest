module xadac
    import xadac_pkg::*;
(
    input logic clk,
    input logic rstn,


);


endmodule
