module xadac_vload_unit
    import xadac_pkg::*;
(
    input logic clk_i,
    input logic rst_ni,

    xadac_ex_if.Slave slv,
    obi_if.Master     obi
);

endmodule
