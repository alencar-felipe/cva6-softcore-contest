module xadac_vactv_unit
    import xadac_ex_if::*;
(
    input logic clk_i,
    input logic rst_ni,

    xadac_ex_if.Slave slv,
    obi_if.Master     obi
);

endmodule
